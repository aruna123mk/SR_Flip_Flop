`include "sr_seqitem.sv"   // Sequence item definition
`include "sr_seq.sv"       // Sequence definition
`include "sr_seqr.sv"      // Sequencer definition
`include "sr_drv.sv"       // Driver definition
`include "sr_mon.sv"       // Monitor definition
`include "sr_agt.sv"       // Agent definition
`include "sr_scbd.sv"      // Scoreboard definition
`include "sr_env.sv"       // Environment definition
`include "sr_test.sv"      // Test definition
